/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:18:22 2023
// Last Modified  : Wed Sep 27 14:18:24 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_slv_env_pkg.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

