/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:08:12 2023
// Last Modified  : Wed Sep 27 14:08:14 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_mas_env_cfg.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

