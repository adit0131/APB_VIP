/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:21:52 2023
// Last Modified  : Wed Sep 27 14:22:28 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_tb_top.sv
// Module Name 	  : 
// Project Name	  : APB_VIP 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

