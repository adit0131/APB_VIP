/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:17:22 2023
// Last Modified  : Wed Sep 27 14:17:23 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_slv_env_cfg.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

