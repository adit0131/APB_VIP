/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:17:43 2023
// Last Modified  : Wed Sep 27 14:17:44 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_slv_sb.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

