/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:09:42 2023
// Last Modified  : Tue Oct  3 14:53:55 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_mas_env_pkg.sv
// Package Name 	: apb_mas_env_pkg 
// Project Name	  : APB_VIP
// Description	  : 
//////////////////////////////////////////////////////////////////////////

`ifndef APB_MAS_ENV_PKG_SV
`define APB_MAS_ENV_PKG_SV 

`include "apb_mas_inf.sv"

package apb_mas_env_pkg;

  import uvm_pkg::*;
 
  `include "uvm_macros.svh";
  
  `include "apb_mas_define.sv";
  `include "apb_mas_agent_cfg.sv";
  `include "apb_mas_seq_item.sv";
  `include "apb_mas_env_cfg.sv";
  `include "apb_mas_drv.sv";
  `include "apb_mas_seqr.sv";
  `include "apb_mas_mon.sv";
  `include "apb_mas_agent.sv";
  `include "apb_mas_base_seqs.sv";
  `include "apb_mas_collector.sv";
  `include "apb_mas_checker.sv";
  `include "apb_mas_sb.sv";  
  `include "apb_mas_env.sv";
 
endpackage

`endif 
