/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:11:55 2023
// Last Modified  : Wed Sep 27 14:11:57 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_mas_sb.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

