/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:05:54 2023
// Last Modified  : Wed Sep 27 14:05:57 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_mas_mon.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

