/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:09:42 2023
// Last Modified  : Wed Sep 27 14:09:44 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_mas_env_pkg.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

