/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:06:18 2023
// Last Modified  : Wed Sep 27 14:06:26 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_mas_agent.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

