/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:05:22 2023
// Last Modified  : Wed Sep 27 14:05:29 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_mas_drv.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

