/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:07:04 2023
// Last Modified  : Wed Sep 27 14:07:05 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_mas_agent_cfg.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

