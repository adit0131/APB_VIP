/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:19:54 2023
// Last Modified  : Wed Sep 27 14:23:09 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_base_test.sv
// Class Name 	  : 
// Project Name	  : APB_VIP 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

