/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:16:55 2023
// Last Modified  : Wed Sep 27 14:16:57 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_slv_env.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

