/////////////////////////////////////////////////////////////////////////
// Company        : SCALEDGE 
// Engineer       : Aditya Mishra 
// Create Date    : Wed Sep 27 14:07:31 2023
// Last Modified  : Wed Sep 27 14:07:47 2023
// Modified By    : Aditya Mishra 
// File Name   	  : apb_mas_env.sv
// Class Name 	  : 
// Project Name	  : 
// Description	  : 
//////////////////////////////////////////////////////////////////////////

